
module __(skeletor-underscore-proj-name)__ #(parameter N=8)
   (
  input	 a,
  output b)
  // TODO
endmodule 
