
module __(skeletor-underscore-proj-name)__ #(parameter N=8)
   (
  input [N-1:0]	 a,
  output [N-1:0] b);
  // TODO
endmodule 
